library ieee;
use ieee.std_logic_1164.all;

package MicDataPkg is

constant MIC_DAT_C : std_logic_vector := (
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0',
'0',
'1',
'0',
'1',
'0',
'1',
'0'
);
end package MicDataPkg;
